`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/06/2024 02:38:12 PM
// Design Name: 
// Module Name: uart_rx
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module uart_rx
    #(
     parameter DBIT = 8,    // data bit
               SB_TICK = 16  // tick for stop bit
    )
    (
     input logic clk, reset,
     input rx, s_tick,
     output logic rx_done_tick,
     output logic [7:0] dout 
    );
    
    // fsm state type
    typedef enum {idle, start, data, stop} state_type;
    
    // signal declaration 
    state_type state_reg, state_next;
    logic [3:0] s_reg, s_next;  // number of tick
    logic [2:0] n_reg, n_next;  // number of data bit
    logic [7:0] b_reg, b_next;  // data (rx  b[7:1])
    
    // FSM
    // state register
    always_ff @(posedge clk, posedge reset)
    begin
        if(reset)
        begin
            state_reg <= idle;
            s_reg <= 0;
            n_reg <= 0;
            b_reg <= 0;
        end
        else
        begin
            state_reg <= state_next;
            s_reg <= s_next;
            n_reg <= n_next;
            b_reg <= b_next;
        end
    end
    
    // next state logic
    always_comb
    begin
        state_next = state_reg;
        rx_done_tick = 0;
        s_next = s_reg;
        n_next = n_reg;
        b_next = b_reg;
        case(state_reg)
        idle:
            if(~rx) // start bit
            begin
                state_next = start;
                s_next = 0;
            end
        start:
            if(s_tick==1)
            begin
                if(s_reg==7)
                begin
                    state_next = data;
                    s_next = 0;
                    n_next = 0;
                end
                else
                    s_next = s_reg + 1;
            end
        data:
        begin
            if(s_tick==1)
            begin
                if(s_reg==15)
                begin
                    s_next = 0;
                    b_next = {rx, b_reg[7:1]};
                    if(n_reg == (DBIT-1))
                    begin
                        state_next = stop;
                    end
                    else
                        n_next = n_reg + 1;
                end
                else
                    s_next = s_reg + 1;
            end
        end
        stop:
        begin
            if(s_tick==1)
            begin
                if(s_reg==(SB_TICK-1))
                begin
                    state_next = idle;
                    rx_done_tick = 1;
                end
                else
                    s_next = s_reg + 1;
            end
        end
        endcase
    end
    
    // output logic 
    assign dout = b_reg;
endmodule
